
//===============================================================================================================================================//
//-----------------------------------------------------------MEM   SEQUENCER---------------------------------------------------------------------//
//===============================================================================================================================================//


class mem_sequencer extends uvm_sequencer#(ethernet_sequence_item);

	`uvm_component_utils(mem_sequencer)


	//===================================== component construction ===================================//

		function  new(string name="mem_sequencer",uvm_component parent);
			super.new(name,parent);
		endfunction
	
	
endclass
